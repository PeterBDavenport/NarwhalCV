module NarshalCV();
	
endmodule 